module next_byte_gen_tb


endmodule