`define next_adr_rom_input_size 9
`define next_adr_rom_output_size 9
module next_adr_rom(input [8:0] data_in, output [8:0] data_out);
        begin
            always@*
            begin
                case(data_in)

					9'b000000000: data_out <= 9'd0;
					9'b000000001: data_out <= 9'd0;
					9'b000000010: data_out <= 9'd0;
					9'b000000011: data_out <= 9'd0;
					9'b000000100: data_out <= 9'd0;
					9'b000000101: data_out <= 9'd0;
					9'b000000110: data_out <= 9'd0;
					9'b000000111: data_out <= 9'd0;
					9'b000001000: data_out <= 9'd0;
					9'b000001001: data_out <= 9'd0;
					9'b000001010: data_out <= 9'd0;
					9'b000001011: data_out <= 9'd268;
					9'b000001100: data_out <= 9'd268;
					9'b000001101: data_out <= 9'd268;
					9'b000001110: data_out <= 9'd269;
					9'b000001111: data_out <= 9'd269;
					9'b000010000: data_out <= 9'd0;
					9'b000010001: data_out <= 9'd0;
					9'b000010010: data_out <= 9'd0;
					9'b000010011: data_out <= 9'd0;
					9'b000010100: data_out <= 9'd0;
					9'b000010101: data_out <= 9'd0;
					9'b000010110: data_out <= 9'd0;
					9'b000010111: data_out <= 9'd275;
					9'b000011000: data_out <= 9'd0;
					9'b000011001: data_out <= 9'd0;
					9'b000011010: data_out <= 9'd0;
					9'b000011011: data_out <= 9'd0;
					9'b000011100: data_out <= 9'd0;
					9'b000011101: data_out <= 9'd0;
					9'b000011110: data_out <= 9'd0;
					9'b000011111: data_out <= 9'd0;
					9'b000100000: data_out <= 9'd0;
					9'b000100001: data_out <= 9'd0;
					9'b000100010: data_out <= 9'd268;
					9'b000100011: data_out <= 9'd268;
					9'b000100100: data_out <= 9'd268;
					9'b000100101: data_out <= 9'd268;
					9'b000100110: data_out <= 9'd0;
					9'b000100111: data_out <= 9'd0;
					9'b000101000: data_out <= 9'd0;
					9'b000101001: data_out <= 9'd0;
					9'b000101010: data_out <= 9'd0;
					9'b000101011: data_out <= 9'd0;
					9'b000101100: data_out <= 9'd0;
					9'b000101101: data_out <= 9'd0;
					9'b000101110: data_out <= 9'd0;
					9'b000101111: data_out <= 9'd0;
					9'b000110000: data_out <= 9'd308;
					9'b000110001: data_out <= 9'd314;
					9'b000110010: data_out <= 9'd0;
					9'b000110011: data_out <= 9'd0;
					9'b000110100: data_out <= 9'd0;
					9'b000110101: data_out <= 9'd0;
					9'b000110110: data_out <= 9'd0;
					9'b000110111: data_out <= 9'd0;
					9'b000111000: data_out <= 9'd0;
					9'b000111001: data_out <= 9'd0;
					9'b000111010: data_out <= 9'd0;
					9'b000111011: data_out <= 9'd0;
					9'b000111100: data_out <= 9'd0;
					9'b000111101: data_out <= 9'd0;
					9'b000111110: data_out <= 9'd0;
					9'b000111111: data_out <= 9'd0;
					9'b001000000: data_out <= 9'd0;
					9'b001000001: data_out <= 9'd0;
					9'b001000010: data_out <= 9'd0;
					9'b001000011: data_out <= 9'd0;
					9'b001000100: data_out <= 9'd0;
					9'b001000101: data_out <= 9'd0;
					9'b001000110: data_out <= 9'd0;
					9'b001000111: data_out <= 9'd0;
					9'b001001000: data_out <= 9'd0;
					9'b001001001: data_out <= 9'd0;
					9'b001001010: data_out <= 9'd0;
					9'b001001011: data_out <= 9'd0;
					9'b001001100: data_out <= 9'd0;
					9'b001001101: data_out <= 9'd0;
					9'b001001110: data_out <= 9'd0;
					9'b001001111: data_out <= 9'd0;
					9'b001010000: data_out <= 9'd0;
					9'b001010001: data_out <= 9'd310;
					9'b001010010: data_out <= 9'd317;
					9'b001010011: data_out <= 9'd0;
					9'b001010100: data_out <= 9'd0;
					9'b001010101: data_out <= 9'd0;
					9'b001010110: data_out <= 9'd0;
					9'b001010111: data_out <= 9'd0;
					9'b001011000: data_out <= 9'd0;
					9'b001011001: data_out <= 9'd256;
					9'b001011010: data_out <= 9'd260;
					9'b001011011: data_out <= 9'd261;
					9'b001011100: data_out <= 9'd258;
					9'b001011101: data_out <= 9'd265;
					9'b001011110: data_out <= 9'd266;
					9'b001011111: data_out <= 9'd263;
					9'b001100000: data_out <= 9'd0;
					9'b001100001: data_out <= 9'd0;
					9'b001100010: data_out <= 9'd272;
					9'b001100011: data_out <= 9'd306;
					9'b001100100: data_out <= 9'd0;
					9'b001100101: data_out <= 9'd0;
					9'b001100110: data_out <= 9'd0;
					9'b001100111: data_out <= 9'd307;
					9'b001101000: data_out <= 9'd0;
					9'b001101001: data_out <= 9'd0;
					9'b001101010: data_out <= 9'd271;
					9'b001101011: data_out <= 9'd0;
					9'b001101100: data_out <= 9'd0;
					9'b001101101: data_out <= 9'd0;
					9'b001101110: data_out <= 9'd270;
					9'b001101111: data_out <= 9'd0;
					9'b001110000: data_out <= 9'd0;
					9'b001110001: data_out <= 9'd0;
					9'b001110010: data_out <= 9'd294;
					9'b001110011: data_out <= 9'd0;
					9'b001110100: data_out <= 9'd0;
					9'b001110101: data_out <= 9'd0;
					9'b001110110: data_out <= 9'd293;
					9'b001110111: data_out <= 9'd0;
					9'b001111000: data_out <= 9'd0;
					9'b001111001: data_out <= 9'd0;
					9'b001111010: data_out <= 9'd0;
					9'b001111011: data_out <= 9'd0;
					9'b001111100: data_out <= 9'd0;
					9'b001111101: data_out <= 9'd0;
					9'b001111110: data_out <= 9'd0;
					9'b001111111: data_out <= 9'd0;
					9'b010000000: data_out <= 9'd0;
					9'b010000001: data_out <= 9'd0;
					9'b010000010: data_out <= 9'd0;
					9'b010000011: data_out <= 9'd0;
					9'b010000100: data_out <= 9'd0;
					9'b010000101: data_out <= 9'd0;
					9'b010000110: data_out <= 9'd0;
					9'b010000111: data_out <= 9'd0;
					9'b010001000: data_out <= 9'd0;
					9'b010001001: data_out <= 9'd0;
					9'b010001010: data_out <= 9'd0;
					9'b010001011: data_out <= 9'd300;
					9'b010001100: data_out <= 9'd302;
					9'b010001101: data_out <= 9'd299;
					9'b010001110: data_out <= 9'd287;
					9'b010001111: data_out <= 9'd288;
					9'b010010000: data_out <= 9'd305;
					9'b010010001: data_out <= 9'd0;
					9'b010010010: data_out <= 9'd0;
					9'b010010011: data_out <= 9'd0;
					9'b010010100: data_out <= 9'd0;
					9'b010010101: data_out <= 9'd278;
					9'b010010110: data_out <= 9'd278;
					9'b010010111: data_out <= 9'd286;
					9'b010011000: data_out <= 9'd286;
					9'b010011001: data_out <= 9'd0;
					9'b010011010: data_out <= 9'd0;
					9'b010011011: data_out <= 9'd0;
					9'b010011100: data_out <= 9'd0;
					9'b010011101: data_out <= 9'd0;
					9'b010011110: data_out <= 9'd0;
					9'b010011111: data_out <= 9'd0;
					9'b010100000: data_out <= 9'd0;
					9'b010100001: data_out <= 9'd0;
					9'b010100010: data_out <= 9'd0;
					9'b010100011: data_out <= 9'd0;
					9'b010100100: data_out <= 9'd0;
					9'b010100101: data_out <= 9'd0;
					9'b010100110: data_out <= 9'd0;
					9'b010100111: data_out <= 9'd0;
					9'b010101000: data_out <= 9'd0;
					9'b010101001: data_out <= 9'd0;
					9'b010101010: data_out <= 9'd0;
					9'b010101011: data_out <= 9'd0;
					9'b010101100: data_out <= 9'd0;
					9'b010101101: data_out <= 9'd0;
					9'b010101110: data_out <= 9'd0;
					9'b010101111: data_out <= 9'd0;
					9'b010110000: data_out <= 9'd0;
					9'b010110001: data_out <= 9'd0;
					9'b010110010: data_out <= 9'd0;
					9'b010110011: data_out <= 9'd0;
					9'b010110100: data_out <= 9'd0;
					9'b010110101: data_out <= 9'd0;
					9'b010110110: data_out <= 9'd0;
					9'b010110111: data_out <= 9'd0;
					9'b010111000: data_out <= 9'd0;
					9'b010111001: data_out <= 9'd0;
					9'b010111010: data_out <= 9'd0;
					9'b010111011: data_out <= 9'd0;
					9'b010111100: data_out <= 9'd0;
					9'b010111101: data_out <= 9'd0;
					9'b010111110: data_out <= 9'd0;
					9'b010111111: data_out <= 9'd0;
					9'b011000000: data_out <= 9'd0;
					9'b011000001: data_out <= 9'd0;
					9'b011000010: data_out <= 9'd0;
					9'b011000011: data_out <= 9'd0;
					9'b011000100: data_out <= 9'd0;
					9'b011000101: data_out <= 9'd0;
					9'b011000110: data_out <= 9'd0;
					9'b011000111: data_out <= 9'd0;
					9'b011001000: data_out <= 9'd0;
					9'b011001001: data_out <= 9'd0;
					9'b011001010: data_out <= 9'd0;
					9'b011001011: data_out <= 9'd0;
					9'b011001100: data_out <= 9'd0;
					9'b011001101: data_out <= 9'd0;
					9'b011001110: data_out <= 9'd0;
					9'b011001111: data_out <= 9'd0;
					9'b011010000: data_out <= 9'd0;
					9'b011010001: data_out <= 9'd0;
					9'b011010010: data_out <= 9'd0;
					9'b011010011: data_out <= 9'd0;
					9'b011010100: data_out <= 9'd0;
					9'b011010101: data_out <= 9'd0;
					9'b011010110: data_out <= 9'd0;
					9'b011010111: data_out <= 9'd0;
					9'b011011000: data_out <= 9'd0;
					9'b011011001: data_out <= 9'd0;
					9'b011011010: data_out <= 9'd0;
					9'b011011011: data_out <= 9'd0;
					9'b011011100: data_out <= 9'd0;
					9'b011011101: data_out <= 9'd0;
					9'b011011110: data_out <= 9'd0;
					9'b011011111: data_out <= 9'd0;
					9'b011100000: data_out <= 9'd0;
					9'b011100001: data_out <= 9'd0;
					9'b011100010: data_out <= 9'd0;
					9'b011100011: data_out <= 9'd0;
					9'b011100100: data_out <= 9'd0;
					9'b011100101: data_out <= 9'd0;
					9'b011100110: data_out <= 9'd0;
					9'b011100111: data_out <= 9'd0;
					9'b011101000: data_out <= 9'd0;
					9'b011101001: data_out <= 9'd0;
					9'b011101010: data_out <= 9'd0;
					9'b011101011: data_out <= 9'd0;
					9'b011101100: data_out <= 9'd0;
					9'b011101101: data_out <= 9'd0;
					9'b011101110: data_out <= 9'd0;
					9'b011101111: data_out <= 9'd0;
					9'b011110000: data_out <= 9'd0;
					9'b011110001: data_out <= 9'd0;
					9'b011110010: data_out <= 9'd0;
					9'b011110011: data_out <= 9'd0;
					9'b011110100: data_out <= 9'd0;
					9'b011110101: data_out <= 9'd0;
					9'b011110110: data_out <= 9'd0;
					9'b011110111: data_out <= 9'd0;
					9'b011111000: data_out <= 9'd0;
					9'b011111001: data_out <= 9'd0;
					9'b011111010: data_out <= 9'd0;
					9'b011111011: data_out <= 9'd0;
					9'b011111100: data_out <= 9'd0;
					9'b011111101: data_out <= 9'd0;
					9'b011111110: data_out <= 9'd0;
					9'b011111111: data_out <= 9'd0;
					9'b100000000: data_out <= 9'd257;
					9'b100000001: data_out <= 9'd0;
					9'b100000010: data_out <= 9'd259;
					9'b100000011: data_out <= 9'd0;
					9'b100000100: data_out <= 9'd259;
					9'b100000101: data_out <= 9'd262;
					9'b100000110: data_out <= 9'd0;
					9'b100000111: data_out <= 9'd264;
					9'b100001000: data_out <= 9'd0;
					9'b100001001: data_out <= 9'd262;
					9'b100001010: data_out <= 9'd267;
					9'b100001011: data_out <= 9'd0;
					9'b100001100: data_out <= 9'd0;
					9'b100001101: data_out <= 9'd0;
					9'b100001110: data_out <= 9'd268;
					9'b100001111: data_out <= 9'd268;
					9'b100010000: data_out <= 9'd273;
					9'b100010001: data_out <= 9'd274;
					9'b100010010: data_out <= 9'd0;
					9'b100010011: data_out <= 9'd276;
					9'b100010100: data_out <= 9'd277;
					9'b100010101: data_out <= 9'd268;
					9'b100010110: data_out <= 9'd279;
					9'b100010111: data_out <= 9'd280;
					9'b100011000: data_out <= 9'd281;
					9'b100011001: data_out <= 9'd282;
					9'b100011010: data_out <= 9'd283;
					9'b100011011: data_out <= 9'd284;
					9'b100011100: data_out <= 9'd285;
					9'b100011101: data_out <= 9'd0;
					9'b100011110: data_out <= 9'd279;
					9'b100011111: data_out <= 9'd268;
					9'b100100000: data_out <= 9'd289;
					9'b100100001: data_out <= 9'd290;
					9'b100100010: data_out <= 9'd291;
					9'b100100011: data_out <= 9'd292;
					9'b100100100: data_out <= 9'd0;
					9'b100100101: data_out <= 9'd268;
					9'b100100110: data_out <= 9'd295;
					9'b100100111: data_out <= 9'd296;
					9'b100101000: data_out <= 9'd297;
					9'b100101001: data_out <= 9'd298;
					9'b100101010: data_out <= 9'd268;
					9'b100101011: data_out <= 9'd269;
					9'b100101100: data_out <= 9'd301;
					9'b100101101: data_out <= 9'd0;
					9'b100101110: data_out <= 9'd303;
					9'b100101111: data_out <= 9'd304;
					9'b100110000: data_out <= 9'd259;
					9'b100110001: data_out <= 9'd268;
					9'b100110010: data_out <= 9'd269;
					9'b100110011: data_out <= 9'd269;
					9'b100110100: data_out <= 9'd309;
					9'b100110101: data_out <= 9'd277;
					9'b100110110: data_out <= 9'd311;
					9'b100110111: data_out <= 9'd312;
					9'b100111000: data_out <= 9'd313;
					9'b100111001: data_out <= 9'd0;
					9'b100111010: data_out <= 9'd315;
					9'b100111011: data_out <= 9'd316;
					9'b100111100: data_out <= 9'd269;
					9'b100111101: data_out <= 9'd318;
					9'b100111110: data_out <= 9'd319;
					9'b100111111: data_out <= 9'd320;
					9'b101000000: data_out <= 9'd0;

                    default: data_out = -1;

                endcase
            end
        end
    endmodule