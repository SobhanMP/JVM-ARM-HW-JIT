`define next_adr_rom_input_size 9
`define next_adr_rom_output_size 9
module next_adr_rom(input [8:0] data_in, output [8:0] data_out);
        begin
            always@*
            begin
                case(data_in)

					9'b000000000 = 9'd0;
					9'b000000001 = 9'd0;
					9'b000000010 = 9'd0;
					9'b000000011 = 9'd0;
					9'b000000100 = 9'd0;
					9'b000000101 = 9'd0;
					9'b000000110 = 9'd0;
					9'b000000111 = 9'd0;
					9'b000001000 = 9'd0;
					9'b000001001 = 9'd0;
					9'b000001010 = 9'd0;
					9'b000001011 = 9'd0;
					9'b000001100 = 9'd0;
					9'b000001101 = 9'd0;
					9'b000001110 = 9'd0;
					9'b000001111 = 9'd0;
					9'b000010000 = 9'd0;
					9'b000010001 = 9'd0;
					9'b000010010 = 9'd0;
					9'b000010011 = 9'd0;
					9'b000010100 = 9'd0;
					9'b000010101 = 9'd0;
					9'b000010110 = 9'd0;
					9'b000010111 = 9'd0;
					9'b000011000 = 9'd0;
					9'b000011001 = 9'd0;
					9'b000011010 = 9'd0;
					9'b000011011 = 9'd0;
					9'b000011100 = 9'd0;
					9'b000011101 = 9'd0;
					9'b000011110 = 9'd0;
					9'b000011111 = 9'd0;
					9'b000100000 = 9'd0;
					9'b000100001 = 9'd0;
					9'b000100010 = 9'd0;
					9'b000100011 = 9'd0;
					9'b000100100 = 9'd0;
					9'b000100101 = 9'd0;
					9'b000100110 = 9'd0;
					9'b000100111 = 9'd0;
					9'b000101000 = 9'd0;
					9'b000101001 = 9'd0;
					9'b000101010 = 9'd0;
					9'b000101011 = 9'd0;
					9'b000101100 = 9'd0;
					9'b000101101 = 9'd0;
					9'b000101110 = 9'd0;
					9'b000101111 = 9'd0;
					9'b000110000 = 9'd0;
					9'b000110001 = 9'd0;
					9'b000110010 = 9'd0;
					9'b000110011 = 9'd0;
					9'b000110100 = 9'd0;
					9'b000110101 = 9'd0;
					9'b000110110 = 9'd0;
					9'b000110111 = 9'd0;
					9'b000111000 = 9'd0;
					9'b000111001 = 9'd0;
					9'b000111010 = 9'd0;
					9'b000111011 = 9'd0;
					9'b000111100 = 9'd0;
					9'b000111101 = 9'd0;
					9'b000111110 = 9'd0;
					9'b000111111 = 9'd0;
					9'b001000000 = 9'd0;
					9'b001000001 = 9'd0;
					9'b001000010 = 9'd0;
					9'b001000011 = 9'd0;
					9'b001000100 = 9'd0;
					9'b001000101 = 9'd0;
					9'b001000110 = 9'd0;
					9'b001000111 = 9'd0;
					9'b001001000 = 9'd0;
					9'b001001001 = 9'd0;
					9'b001001010 = 9'd0;
					9'b001001011 = 9'd0;
					9'b001001100 = 9'd0;
					9'b001001101 = 9'd0;
					9'b001001110 = 9'd0;
					9'b001001111 = 9'd0;
					9'b001010000 = 9'd0;
					9'b001010001 = 9'd0;
					9'b001010010 = 9'd0;
					9'b001010011 = 9'd0;
					9'b001010100 = 9'd0;
					9'b001010101 = 9'd0;
					9'b001010110 = 9'd0;
					9'b001010111 = 9'd0;
					9'b001011000 = 9'd0;
					9'b001011001 = 9'd0;
					9'b001011010 = 9'd0;
					9'b001011011 = 9'd0;
					9'b001011100 = 9'd0;
					9'b001011101 = 9'd0;
					9'b001011110 = 9'd0;
					9'b001011111 = 9'd0;
					9'b001100000 = 9'd256;
					9'b001100001 = 9'd0;
					9'b001100010 = 9'd0;
					9'b001100011 = 9'd0;
					9'b001100100 = 9'd258;
					9'b001100101 = 9'd0;
					9'b001100110 = 9'd0;
					9'b001100111 = 9'd0;
					9'b001101000 = 9'd0;
					9'b001101001 = 9'd0;
					9'b001101010 = 9'd0;
					9'b001101011 = 9'd0;
					9'b001101100 = 9'd0;
					9'b001101101 = 9'd0;
					9'b001101110 = 9'd0;
					9'b001101111 = 9'd0;
					9'b001110000 = 9'd0;
					9'b001110001 = 9'd0;
					9'b001110010 = 9'd0;
					9'b001110011 = 9'd0;
					9'b001110100 = 9'd0;
					9'b001110101 = 9'd0;
					9'b001110110 = 9'd0;
					9'b001110111 = 9'd0;
					9'b001111000 = 9'd0;
					9'b001111001 = 9'd0;
					9'b001111010 = 9'd0;
					9'b001111011 = 9'd0;
					9'b001111100 = 9'd0;
					9'b001111101 = 9'd0;
					9'b001111110 = 9'd0;
					9'b001111111 = 9'd0;
					9'b010000000 = 9'd0;
					9'b010000001 = 9'd0;
					9'b010000010 = 9'd0;
					9'b010000011 = 9'd0;
					9'b010000100 = 9'd0;
					9'b010000101 = 9'd0;
					9'b010000110 = 9'd0;
					9'b010000111 = 9'd0;
					9'b010001000 = 9'd0;
					9'b010001001 = 9'd0;
					9'b010001010 = 9'd0;
					9'b010001011 = 9'd0;
					9'b010001100 = 9'd0;
					9'b010001101 = 9'd0;
					9'b010001110 = 9'd0;
					9'b010001111 = 9'd0;
					9'b010010000 = 9'd0;
					9'b010010001 = 9'd0;
					9'b010010010 = 9'd0;
					9'b010010011 = 9'd0;
					9'b010010100 = 9'd0;
					9'b010010101 = 9'd0;
					9'b010010110 = 9'd0;
					9'b010010111 = 9'd0;
					9'b010011000 = 9'd0;
					9'b010011001 = 9'd0;
					9'b010011010 = 9'd0;
					9'b010011011 = 9'd0;
					9'b010011100 = 9'd0;
					9'b010011101 = 9'd0;
					9'b010011110 = 9'd0;
					9'b010011111 = 9'd0;
					9'b010100000 = 9'd0;
					9'b010100001 = 9'd0;
					9'b010100010 = 9'd0;
					9'b010100011 = 9'd0;
					9'b010100100 = 9'd0;
					9'b010100101 = 9'd0;
					9'b010100110 = 9'd0;
					9'b010100111 = 9'd0;
					9'b010101000 = 9'd0;
					9'b010101001 = 9'd0;
					9'b010101010 = 9'd0;
					9'b010101011 = 9'd0;
					9'b010101100 = 9'd0;
					9'b010101101 = 9'd0;
					9'b010101110 = 9'd0;
					9'b010101111 = 9'd0;
					9'b010110000 = 9'd0;
					9'b010110001 = 9'd0;
					9'b010110010 = 9'd0;
					9'b010110011 = 9'd0;
					9'b010110100 = 9'd0;
					9'b010110101 = 9'd0;
					9'b010110110 = 9'd0;
					9'b010110111 = 9'd0;
					9'b010111000 = 9'd0;
					9'b010111001 = 9'd0;
					9'b010111010 = 9'd0;
					9'b010111011 = 9'd0;
					9'b010111100 = 9'd0;
					9'b010111101 = 9'd0;
					9'b010111110 = 9'd0;
					9'b010111111 = 9'd0;
					9'b011000000 = 9'd0;
					9'b011000001 = 9'd0;
					9'b011000010 = 9'd0;
					9'b011000011 = 9'd0;
					9'b011000100 = 9'd0;
					9'b011000101 = 9'd0;
					9'b011000110 = 9'd0;
					9'b011000111 = 9'd0;
					9'b011001000 = 9'd0;
					9'b011001001 = 9'd0;
					9'b011001010 = 9'd0;
					9'b011001011 = 9'd0;
					9'b011001100 = 9'd0;
					9'b011001101 = 9'd0;
					9'b011001110 = 9'd0;
					9'b011001111 = 9'd0;
					9'b011010000 = 9'd0;
					9'b011010001 = 9'd0;
					9'b011010010 = 9'd0;
					9'b011010011 = 9'd0;
					9'b011010100 = 9'd0;
					9'b011010101 = 9'd0;
					9'b011010110 = 9'd0;
					9'b011010111 = 9'd0;
					9'b011011000 = 9'd0;
					9'b011011001 = 9'd0;
					9'b011011010 = 9'd0;
					9'b011011011 = 9'd0;
					9'b011011100 = 9'd0;
					9'b011011101 = 9'd0;
					9'b011011110 = 9'd0;
					9'b011011111 = 9'd0;
					9'b011100000 = 9'd0;
					9'b011100001 = 9'd0;
					9'b011100010 = 9'd0;
					9'b011100011 = 9'd0;
					9'b011100100 = 9'd0;
					9'b011100101 = 9'd0;
					9'b011100110 = 9'd0;
					9'b011100111 = 9'd0;
					9'b011101000 = 9'd0;
					9'b011101001 = 9'd0;
					9'b011101010 = 9'd0;
					9'b011101011 = 9'd0;
					9'b011101100 = 9'd0;
					9'b011101101 = 9'd0;
					9'b011101110 = 9'd0;
					9'b011101111 = 9'd0;
					9'b011110000 = 9'd0;
					9'b011110001 = 9'd0;
					9'b011110010 = 9'd0;
					9'b011110011 = 9'd0;
					9'b011110100 = 9'd0;
					9'b011110101 = 9'd0;
					9'b011110110 = 9'd0;
					9'b011110111 = 9'd0;
					9'b011111000 = 9'd0;
					9'b011111001 = 9'd0;
					9'b011111010 = 9'd0;
					9'b011111011 = 9'd0;
					9'b011111100 = 9'd0;
					9'b011111101 = 9'd0;
					9'b011111110 = 9'd0;
					9'b011111111 = 9'd0;
					9'b100000000 = 9'd257;
					9'b100000001 = 9'd0;
					9'b100000010 = 9'd257;

                    default: data_out = -1;

                endcase
            end
        end
    endmodule