// input: opcode of jvm instruction
// output: number of bytes after that instruction
module count_rom(output reg[4:0] count, input wire [7:0] opcode);
    always @(opcode) begin
        case (address) 
            8'b0000000: count = 5'd0;
            8'b0000000: count = 5'd0;
            8'b0000001: count = 5'd0;
            8'b0000001: count = 5'd0;
            8'b0000010: count = 5'd0;
            8'b0000010: count = 5'd0;
            8'b0000011: count = 5'd0;
            8'b0000011: count = 5'd0;
            8'b0000100: count = 5'd0;
            8'b0000100: count = 5'd0;
            8'b0000101: count = 5'd0;
            8'b0000101: count = 5'd0;
            8'b0000110: count = 5'd0;
            8'b0000110: count = 5'd0;
            8'b0000111: count = 5'd0;
            8'b0000111: count = 5'd0;
            8'b0001000: count = 5'd1;
            8'b0001000: count = 5'd2;
            8'b0001001: count = 5'd1;
            8'b0001001: count = 5'd2;
            8'b0001010: count = 5'd2;
            8'b0001010: count = 5'd1;
            8'b0001011: count = 5'd1;
            8'b0001011: count = 5'd1;
            8'b0001100: count = 5'd1;
            8'b0001100: count = 5'd1;
            8'b0001101: count = 5'd0;
            8'b0001101: count = 5'd0;
            8'b0001110: count = 5'd0;
            8'b0001110: count = 5'd0;
            8'b0001111: count = 5'd0;
            8'b0001111: count = 5'd0;
            8'b0010000: count = 5'd0;
            8'b0010000: count = 5'd0;
            8'b0010001: count = 5'd0;
            8'b0010001: count = 5'd0;
            8'b0010010: count = 5'd0;
            8'b0010010: count = 5'd0;
            8'b0010011: count = 5'd0;
            8'b0010011: count = 5'd0;
            8'b0010100: count = 5'd0;
            8'b0010100: count = 5'd0;
            8'b0010101: count = 5'd0;
            8'b0010101: count = 5'd0;
            8'b0010110: count = 5'd0;
            8'b0010110: count = 5'd0;
            8'b0010111: count = 5'd0;
            8'b0010111: count = 5'd0;
            8'b0011000: count = 5'd0;
            8'b0011000: count = 5'd0;
            8'b0011001: count = 5'd0;
            8'b0011001: count = 5'd0;
            8'b0011010: count = 5'd0;
            8'b0011010: count = 5'd0;
            8'b0011011: count = 5'd1;
            8'b0011011: count = 5'd1;
            8'b0011100: count = 5'd1;
            8'b0011100: count = 5'd1;
            8'b0011101: count = 5'd1;
            8'b0011101: count = 5'd0;
            8'b0011110: count = 5'd0;
            8'b0011110: count = 5'd0;
            8'b0011111: count = 5'd0;
            8'b0011111: count = 5'd0;
            8'b0100000: count = 5'd0;
            8'b0100000: count = 5'd0;
            8'b0100001: count = 5'd0;
            8'b0100001: count = 5'd0;
            8'b0100010: count = 5'd0;
            8'b0100010: count = 5'd0;
            8'b0100011: count = 5'd0;
            8'b0100011: count = 5'd0;
            8'b0100100: count = 5'd0;
            8'b0100100: count = 5'd0;
            8'b0100101: count = 5'd0;
            8'b0100101: count = 5'd0;
            8'b0100110: count = 5'd0;
            8'b0100110: count = 5'd0;
            8'b0100111: count = 5'd0;
            8'b0100111: count = 5'd0;
            8'b0101000: count = 5'd0;
            8'b0101000: count = 5'd0;
            8'b0101001: count = 5'd0;
            8'b0101001: count = 5'd0;
            8'b0101010: count = 5'd0;
            8'b0101010: count = 5'd0;
            8'b0101011: count = 5'd0;
            8'b0101011: count = 5'd0;
            8'b0101100: count = 5'd0;
            8'b0101100: count = 5'd0;
            8'b0101101: count = 5'd0;
            8'b0101101: count = 5'd0;
            8'b0101110: count = 5'd0;
            8'b0101110: count = 5'd0;
            8'b0101111: count = 5'd0;
            8'b0101111: count = 5'd0;
            8'b0110000: count = 5'd0;
            8'b0110000: count = 5'd0;
            8'b0110001: count = 5'd0;
            8'b0110001: count = 5'd0;
            8'b0110010: count = 5'd0;
            8'b0110010: count = 5'd0;
            8'b0110011: count = 5'd0;
            8'b0110011: count = 5'd0;
            8'b0110100: count = 5'd0;
            8'b0110100: count = 5'd0;
            8'b0110101: count = 5'd0;
            8'b0110101: count = 5'd0;
            8'b0110110: count = 5'd0;
            8'b0110110: count = 5'd0;
            8'b0110111: count = 5'd0;
            8'b0110111: count = 5'd0;
            8'b0111000: count = 5'd0;
            8'b0111000: count = 5'd0;
            8'b0111001: count = 5'd0;
            8'b0111001: count = 5'd0;
            8'b0111010: count = 5'd0;
            8'b0111010: count = 5'd0;
            8'b0111011: count = 5'd0;
            8'b0111011: count = 5'd0;
            8'b0111100: count = 5'd0;
            8'b0111100: count = 5'd0;
            8'b0111101: count = 5'd0;
            8'b0111101: count = 5'd0;
            8'b0111110: count = 5'd0;
            8'b0111110: count = 5'd0;
            8'b0111111: count = 5'd0;
            8'b0111111: count = 5'd0;
            8'b1000000: count = 5'd0;
            8'b1000000: count = 5'd0;
            8'b1000001: count = 5'd0;
            8'b1000001: count = 5'd0;
            8'b1000010: count = 5'd2;
            8'b1000010: count = 5'd0;
            8'b1000011: count = 5'd0;
            8'b1000011: count = 5'd0;
            8'b1000100: count = 5'd0;
            8'b1000100: count = 5'd0;
            8'b1000101: count = 5'd0;
            8'b1000101: count = 5'd0;
            8'b1000110: count = 5'd0;
            8'b1000110: count = 5'd0;
            8'b1000111: count = 5'd0;
            8'b1000111: count = 5'd0;
            8'b1001000: count = 5'd0;
            8'b1001000: count = 5'd0;
            8'b1001001: count = 5'd0;
            8'b1001001: count = 5'd0;
            8'b1001010: count = 5'd0;
            8'b1001010: count = 5'd0;
            8'b1001011: count = 5'd0;
            8'b1001011: count = 5'd0;
            8'b1001100: count = 5'd0;
            8'b1001100: count = 5'd2;
            8'b1001101: count = 5'd2;
            8'b1001101: count = 5'd2;
            8'b1001110: count = 5'd2;
            8'b1001110: count = 5'd2;
            8'b1001111: count = 5'd2;
            8'b1001111: count = 5'd2;
            8'b1010000: count = 5'd2;
            8'b1010000: count = 5'd2;
            8'b1010001: count = 5'd2;
            8'b1010001: count = 5'd2;
            8'b1010010: count = 5'd2;
            8'b1010010: count = 5'd2;
            8'b1010011: count = 5'd2;
            8'b1010011: count = 5'd2;
            8'b1010100: count = 5'd2;
            8'b1010100: count = 5'd1;
            8'b1010101: count = 5'd16;
            8'b1010101: count = 5'd8;
            8'b1010110: count = 5'd0;
            8'b1010110: count = 5'd0;
            8'b1010111: count = 5'd0;
            8'b1010111: count = 5'd0;
            8'b1011000: count = 5'd0;
            8'b1011000: count = 5'd0;
            8'b1011001: count = 5'd2;
            8'b1011001: count = 5'd2;
            8'b1011010: count = 5'd2;
            8'b1011010: count = 5'd2;
            8'b1011011: count = 5'd2;
            8'b1011011: count = 5'd2;
            8'b1011100: count = 5'd2;
            8'b1011100: count = 5'd4;
            8'b1011101: count = 5'd4;
            8'b1011101: count = 5'd2;
            8'b1011110: count = 5'd1;
            8'b1011110: count = 5'd2;
            8'b1011111: count = 5'd0;
            8'b1011111: count = 5'd0;
            8'b1100000: count = 5'd2;
            8'b1100000: count = 5'd2;
            8'b1100001: count = 5'd0;
            8'b1100001: count = 5'd0;
            8'b1100010: count = 5'd3;
            8'b1100010: count = 5'd3;
            8'b1100011: count = 5'd2;
            8'b1100011: count = 5'd2;
            8'b1100100: count = 5'd4;
            8'b1100100: count = 5'd4;
            8'b1100101: count = 5'd0;
            8'b1111111: count = 5'd0;
            8'b1111111: count = 5'd0;
            default: count = 5'd0;
        endcase
    end
endmodule