`define inst_adr_rom_input_size 9
`define inst_adr_rom_output_size 3
module inst_adr_rom(input [8:0] data_in, output [2:0] data_out);
        begin
            always@*
            begin
                case(data_in)

					9'b000000000 = 3'd0;
					9'b000000001 = 3'd0;
					9'b000000010 = 3'd0;
					9'b000000011 = 3'd0;
					9'b000000100 = 3'd0;
					9'b000000101 = 3'd0;
					9'b000000110 = 3'd0;
					9'b000000111 = 3'd0;
					9'b000001000 = 3'd0;
					9'b000001001 = 3'd0;
					9'b000001010 = 3'd0;
					9'b000001011 = 3'd0;
					9'b000001100 = 3'd0;
					9'b000001101 = 3'd0;
					9'b000001110 = 3'd0;
					9'b000001111 = 3'd0;
					9'b000010000 = 3'd0;
					9'b000010001 = 3'd0;
					9'b000010010 = 3'd0;
					9'b000010011 = 3'd0;
					9'b000010100 = 3'd0;
					9'b000010101 = 3'd0;
					9'b000010110 = 3'd0;
					9'b000010111 = 3'd0;
					9'b000011000 = 3'd0;
					9'b000011001 = 3'd0;
					9'b000011010 = 3'd0;
					9'b000011011 = 3'd0;
					9'b000011100 = 3'd0;
					9'b000011101 = 3'd0;
					9'b000011110 = 3'd0;
					9'b000011111 = 3'd0;
					9'b000100000 = 3'd0;
					9'b000100001 = 3'd0;
					9'b000100010 = 3'd0;
					9'b000100011 = 3'd0;
					9'b000100100 = 3'd0;
					9'b000100101 = 3'd0;
					9'b000100110 = 3'd0;
					9'b000100111 = 3'd0;
					9'b000101000 = 3'd0;
					9'b000101001 = 3'd0;
					9'b000101010 = 3'd0;
					9'b000101011 = 3'd0;
					9'b000101100 = 3'd0;
					9'b000101101 = 3'd0;
					9'b000101110 = 3'd0;
					9'b000101111 = 3'd0;
					9'b000110000 = 3'd0;
					9'b000110001 = 3'd0;
					9'b000110010 = 3'd0;
					9'b000110011 = 3'd0;
					9'b000110100 = 3'd0;
					9'b000110101 = 3'd0;
					9'b000110110 = 3'd0;
					9'b000110111 = 3'd0;
					9'b000111000 = 3'd0;
					9'b000111001 = 3'd0;
					9'b000111010 = 3'd0;
					9'b000111011 = 3'd0;
					9'b000111100 = 3'd0;
					9'b000111101 = 3'd0;
					9'b000111110 = 3'd0;
					9'b000111111 = 3'd0;
					9'b001000000 = 3'd0;
					9'b001000001 = 3'd0;
					9'b001000010 = 3'd0;
					9'b001000011 = 3'd0;
					9'b001000100 = 3'd0;
					9'b001000101 = 3'd0;
					9'b001000110 = 3'd0;
					9'b001000111 = 3'd0;
					9'b001001000 = 3'd0;
					9'b001001001 = 3'd0;
					9'b001001010 = 3'd0;
					9'b001001011 = 3'd0;
					9'b001001100 = 3'd0;
					9'b001001101 = 3'd0;
					9'b001001110 = 3'd0;
					9'b001001111 = 3'd0;
					9'b001010000 = 3'd0;
					9'b001010001 = 3'd0;
					9'b001010010 = 3'd0;
					9'b001010011 = 3'd0;
					9'b001010100 = 3'd0;
					9'b001010101 = 3'd0;
					9'b001010110 = 3'd0;
					9'b001010111 = 3'd0;
					9'b001011000 = 3'd0;
					9'b001011001 = 3'd0;
					9'b001011010 = 3'd0;
					9'b001011011 = 3'd0;
					9'b001011100 = 3'd0;
					9'b001011101 = 3'd0;
					9'b001011110 = 3'd0;
					9'b001011111 = 3'd0;
					9'b001100000 = 3'd0;
					9'b001100001 = 3'd0;
					9'b001100010 = 3'd0;
					9'b001100011 = 3'd0;
					9'b001100100 = 3'd0;
					9'b001100101 = 3'd0;
					9'b001100110 = 3'd0;
					9'b001100111 = 3'd0;
					9'b001101000 = 3'd0;
					9'b001101001 = 3'd0;
					9'b001101010 = 3'd0;
					9'b001101011 = 3'd0;
					9'b001101100 = 3'd0;
					9'b001101101 = 3'd0;
					9'b001101110 = 3'd0;
					9'b001101111 = 3'd0;
					9'b001110000 = 3'd0;
					9'b001110001 = 3'd0;
					9'b001110010 = 3'd0;
					9'b001110011 = 3'd0;
					9'b001110100 = 3'd0;
					9'b001110101 = 3'd0;
					9'b001110110 = 3'd0;
					9'b001110111 = 3'd0;
					9'b001111000 = 3'd0;
					9'b001111001 = 3'd0;
					9'b001111010 = 3'd0;
					9'b001111011 = 3'd0;
					9'b001111100 = 3'd0;
					9'b001111101 = 3'd0;
					9'b001111110 = 3'd0;
					9'b001111111 = 3'd0;
					9'b010000000 = 3'd0;
					9'b010000001 = 3'd0;
					9'b010000010 = 3'd0;
					9'b010000011 = 3'd0;
					9'b010000100 = 3'd0;
					9'b010000101 = 3'd0;
					9'b010000110 = 3'd0;
					9'b010000111 = 3'd0;
					9'b010001000 = 3'd0;
					9'b010001001 = 3'd0;
					9'b010001010 = 3'd0;
					9'b010001011 = 3'd0;
					9'b010001100 = 3'd0;
					9'b010001101 = 3'd0;
					9'b010001110 = 3'd0;
					9'b010001111 = 3'd0;
					9'b010010000 = 3'd0;
					9'b010010001 = 3'd0;
					9'b010010010 = 3'd0;
					9'b010010011 = 3'd0;
					9'b010010100 = 3'd0;
					9'b010010101 = 3'd0;
					9'b010010110 = 3'd0;
					9'b010010111 = 3'd0;
					9'b010011000 = 3'd0;
					9'b010011001 = 3'd0;
					9'b010011010 = 3'd0;
					9'b010011011 = 3'd0;
					9'b010011100 = 3'd0;
					9'b010011101 = 3'd0;
					9'b010011110 = 3'd0;
					9'b010011111 = 3'd0;
					9'b010100000 = 3'd0;
					9'b010100001 = 3'd0;
					9'b010100010 = 3'd0;
					9'b010100011 = 3'd0;
					9'b010100100 = 3'd0;
					9'b010100101 = 3'd0;
					9'b010100110 = 3'd0;
					9'b010100111 = 3'd0;
					9'b010101000 = 3'd0;
					9'b010101001 = 3'd0;
					9'b010101010 = 3'd0;
					9'b010101011 = 3'd0;
					9'b010101100 = 3'd0;
					9'b010101101 = 3'd0;
					9'b010101110 = 3'd0;
					9'b010101111 = 3'd0;
					9'b010110000 = 3'd0;
					9'b010110001 = 3'd0;
					9'b010110010 = 3'd0;
					9'b010110011 = 3'd0;
					9'b010110100 = 3'd0;
					9'b010110101 = 3'd0;
					9'b010110110 = 3'd0;
					9'b010110111 = 3'd0;
					9'b010111000 = 3'd0;
					9'b010111001 = 3'd0;
					9'b010111010 = 3'd0;
					9'b010111011 = 3'd0;
					9'b010111100 = 3'd0;
					9'b010111101 = 3'd0;
					9'b010111110 = 3'd0;
					9'b010111111 = 3'd0;
					9'b011000000 = 3'd0;
					9'b011000001 = 3'd0;
					9'b011000010 = 3'd0;
					9'b011000011 = 3'd0;
					9'b011000100 = 3'd0;
					9'b011000101 = 3'd0;
					9'b011000110 = 3'd0;
					9'b011000111 = 3'd0;
					9'b011001000 = 3'd0;
					9'b011001001 = 3'd0;
					9'b011001010 = 3'd0;
					9'b011001011 = 3'd0;
					9'b011001100 = 3'd0;
					9'b011001101 = 3'd0;
					9'b011001110 = 3'd0;
					9'b011001111 = 3'd0;
					9'b011010000 = 3'd0;
					9'b011010001 = 3'd0;
					9'b011010010 = 3'd0;
					9'b011010011 = 3'd0;
					9'b011010100 = 3'd0;
					9'b011010101 = 3'd0;
					9'b011010110 = 3'd0;
					9'b011010111 = 3'd0;
					9'b011011000 = 3'd0;
					9'b011011001 = 3'd0;
					9'b011011010 = 3'd0;
					9'b011011011 = 3'd0;
					9'b011011100 = 3'd0;
					9'b011011101 = 3'd0;
					9'b011011110 = 3'd0;
					9'b011011111 = 3'd0;
					9'b011100000 = 3'd0;
					9'b011100001 = 3'd0;
					9'b011100010 = 3'd0;
					9'b011100011 = 3'd0;
					9'b011100100 = 3'd0;
					9'b011100101 = 3'd0;
					9'b011100110 = 3'd0;
					9'b011100111 = 3'd0;
					9'b011101000 = 3'd0;
					9'b011101001 = 3'd0;
					9'b011101010 = 3'd0;
					9'b011101011 = 3'd0;
					9'b011101100 = 3'd0;
					9'b011101101 = 3'd0;
					9'b011101110 = 3'd0;
					9'b011101111 = 3'd0;
					9'b011110000 = 3'd0;
					9'b011110001 = 3'd0;
					9'b011110010 = 3'd0;
					9'b011110011 = 3'd0;
					9'b011110100 = 3'd0;
					9'b011110101 = 3'd0;
					9'b011110110 = 3'd0;
					9'b011110111 = 3'd0;
					9'b011111000 = 3'd0;
					9'b011111001 = 3'd0;
					9'b011111010 = 3'd0;
					9'b011111011 = 3'd0;
					9'b011111100 = 3'd0;
					9'b011111101 = 3'd0;
					9'b011111110 = 3'd0;
					9'b011111111 = 3'd0;
					9'b100000000 = 3'd1;
					9'b100000001 = 3'd2;
					9'b100000010 = 3'd3;

                    default: data_out = -1;

                endcase
            end
        end
    endmodule