`define inst_adr_rom_input_size 9
`define inst_adr_rom_output_size 7
module inst_adr_rom(input [8:0] data_in, output reg [6:0] data_out);
        
            always@*
            begin
                case(data_in)

					9'b000000000: data_out <= 7'd0;
					9'b000000001: data_out <= 7'd0;
					9'b000000010: data_out <= 7'd0;
					9'b000000011: data_out <= 7'd0;
					9'b000000100: data_out <= 7'd0;
					9'b000000101: data_out <= 7'd0;
					9'b000000110: data_out <= 7'd0;
					9'b000000111: data_out <= 7'd0;
					9'b000001000: data_out <= 7'd0;
					9'b000001001: data_out <= 7'd0;
					9'b000001010: data_out <= 7'd0;
					9'b000001011: data_out <= 7'd11;
					9'b000001100: data_out <= 7'd13;
					9'b000001101: data_out <= 7'd14;
					9'b000001110: data_out <= 7'd15;
					9'b000001111: data_out <= 7'd17;
					9'b000010000: data_out <= 7'd0;
					9'b000010001: data_out <= 7'd0;
					9'b000010010: data_out <= 7'd0;
					9'b000010011: data_out <= 7'd0;
					9'b000010100: data_out <= 7'd0;
					9'b000010101: data_out <= 7'd0;
					9'b000010110: data_out <= 7'd0;
					9'b000010111: data_out <= 7'd1;
					9'b000011000: data_out <= 7'd0;
					9'b000011001: data_out <= 7'd0;
					9'b000011010: data_out <= 7'd0;
					9'b000011011: data_out <= 7'd0;
					9'b000011100: data_out <= 7'd0;
					9'b000011101: data_out <= 7'd0;
					9'b000011110: data_out <= 7'd0;
					9'b000011111: data_out <= 7'd0;
					9'b000100000: data_out <= 7'd0;
					9'b000100001: data_out <= 7'd0;
					9'b000100010: data_out <= 7'd26;
					9'b000100011: data_out <= 7'd27;
					9'b000100100: data_out <= 7'd28;
					9'b000100101: data_out <= 7'd29;
					9'b000100110: data_out <= 7'd0;
					9'b000100111: data_out <= 7'd0;
					9'b000101000: data_out <= 7'd0;
					9'b000101001: data_out <= 7'd0;
					9'b000101010: data_out <= 7'd0;
					9'b000101011: data_out <= 7'd0;
					9'b000101100: data_out <= 7'd0;
					9'b000101101: data_out <= 7'd0;
					9'b000101110: data_out <= 7'd0;
					9'b000101111: data_out <= 7'd0;
					9'b000110000: data_out <= 7'd3;
					9'b000110001: data_out <= 7'd3;
					9'b000110010: data_out <= 7'd0;
					9'b000110011: data_out <= 7'd0;
					9'b000110100: data_out <= 7'd0;
					9'b000110101: data_out <= 7'd0;
					9'b000110110: data_out <= 7'd0;
					9'b000110111: data_out <= 7'd0;
					9'b000111000: data_out <= 7'd0;
					9'b000111001: data_out <= 7'd0;
					9'b000111010: data_out <= 7'd0;
					9'b000111011: data_out <= 7'd0;
					9'b000111100: data_out <= 7'd0;
					9'b000111101: data_out <= 7'd0;
					9'b000111110: data_out <= 7'd0;
					9'b000111111: data_out <= 7'd0;
					9'b001000000: data_out <= 7'd0;
					9'b001000001: data_out <= 7'd0;
					9'b001000010: data_out <= 7'd0;
					9'b001000011: data_out <= 7'd0;
					9'b001000100: data_out <= 7'd0;
					9'b001000101: data_out <= 7'd0;
					9'b001000110: data_out <= 7'd0;
					9'b001000111: data_out <= 7'd0;
					9'b001001000: data_out <= 7'd0;
					9'b001001001: data_out <= 7'd0;
					9'b001001010: data_out <= 7'd0;
					9'b001001011: data_out <= 7'd0;
					9'b001001100: data_out <= 7'd0;
					9'b001001101: data_out <= 7'd0;
					9'b001001110: data_out <= 7'd0;
					9'b001001111: data_out <= 7'd0;
					9'b001010000: data_out <= 7'd0;
					9'b001010001: data_out <= 7'd47;
					9'b001010010: data_out <= 7'd40;
					9'b001010011: data_out <= 7'd0;
					9'b001010100: data_out <= 7'd0;
					9'b001010101: data_out <= 7'd0;
					9'b001010110: data_out <= 7'd0;
					9'b001010111: data_out <= 7'd1;
					9'b001011000: data_out <= 7'd3;
					9'b001011001: data_out <= 7'd1;
					9'b001011010: data_out <= 7'd3;
					9'b001011011: data_out <= 7'd5;
					9'b001011100: data_out <= 7'd3;
					9'b001011101: data_out <= 7'd5;
					9'b001011110: data_out <= 7'd9;
					9'b001011111: data_out <= 7'd3;
					9'b001100000: data_out <= 7'd0;
					9'b001100001: data_out <= 7'd0;
					9'b001100010: data_out <= 7'd18;
					9'b001100011: data_out <= 7'd38;
					9'b001100100: data_out <= 7'd0;
					9'b001100101: data_out <= 7'd0;
					9'b001100110: data_out <= 7'd0;
					9'b001100111: data_out <= 7'd38;
					9'b001101000: data_out <= 7'd0;
					9'b001101001: data_out <= 7'd0;
					9'b001101010: data_out <= 7'd18;
					9'b001101011: data_out <= 7'd0;
					9'b001101100: data_out <= 7'd0;
					9'b001101101: data_out <= 7'd0;
					9'b001101110: data_out <= 7'd18;
					9'b001101111: data_out <= 7'd0;
					9'b001110000: data_out <= 7'd0;
					9'b001110001: data_out <= 7'd0;
					9'b001110010: data_out <= 7'd18;
					9'b001110011: data_out <= 7'd0;
					9'b001110100: data_out <= 7'd0;
					9'b001110101: data_out <= 7'd0;
					9'b001110110: data_out <= 7'd47;
					9'b001110111: data_out <= 7'd0;
					9'b001111000: data_out <= 7'd0;
					9'b001111001: data_out <= 7'd0;
					9'b001111010: data_out <= 7'd0;
					9'b001111011: data_out <= 7'd0;
					9'b001111100: data_out <= 7'd0;
					9'b001111101: data_out <= 7'd0;
					9'b001111110: data_out <= 7'd0;
					9'b001111111: data_out <= 7'd0;
					9'b010000000: data_out <= 7'd0;
					9'b010000001: data_out <= 7'd0;
					9'b010000010: data_out <= 7'd0;
					9'b010000011: data_out <= 7'd0;
					9'b010000100: data_out <= 7'd0;
					9'b010000101: data_out <= 7'd0;
					9'b010000110: data_out <= 7'd0;
					9'b010000111: data_out <= 7'd0;
					9'b010001000: data_out <= 7'd0;
					9'b010001001: data_out <= 7'd0;
					9'b010001010: data_out <= 7'd0;
					9'b010001011: data_out <= 7'd47;
					9'b010001100: data_out <= 7'd1;
					9'b010001101: data_out <= 7'd47;
					9'b010001110: data_out <= 7'd40;
					9'b010001111: data_out <= 7'd40;
					9'b010010000: data_out <= 7'd57;
					9'b010010001: data_out <= 7'd0;
					9'b010010010: data_out <= 7'd0;
					9'b010010011: data_out <= 7'd0;
					9'b010010100: data_out <= 7'd0;
					9'b010010101: data_out <= 7'd18;
					9'b010010110: data_out <= 7'd18;
					9'b010010111: data_out <= 7'd38;
					9'b010011000: data_out <= 7'd38;
					9'b010011001: data_out <= 7'd0;
					9'b010011010: data_out <= 7'd0;
					9'b010011011: data_out <= 7'd0;
					9'b010011100: data_out <= 7'd0;
					9'b010011101: data_out <= 7'd0;
					9'b010011110: data_out <= 7'd0;
					9'b010011111: data_out <= 7'd0;
					9'b010100000: data_out <= 7'd0;
					9'b010100001: data_out <= 7'd0;
					9'b010100010: data_out <= 7'd0;
					9'b010100011: data_out <= 7'd0;
					9'b010100100: data_out <= 7'd0;
					9'b010100101: data_out <= 7'd0;
					9'b010100110: data_out <= 7'd0;
					9'b010100111: data_out <= 7'd0;
					9'b010101000: data_out <= 7'd0;
					9'b010101001: data_out <= 7'd0;
					9'b010101010: data_out <= 7'd0;
					9'b010101011: data_out <= 7'd0;
					9'b010101100: data_out <= 7'd0;
					9'b010101101: data_out <= 7'd0;
					9'b010101110: data_out <= 7'd0;
					9'b010101111: data_out <= 7'd0;
					9'b010110000: data_out <= 7'd0;
					9'b010110001: data_out <= 7'd0;
					9'b010110010: data_out <= 7'd0;
					9'b010110011: data_out <= 7'd0;
					9'b010110100: data_out <= 7'd0;
					9'b010110101: data_out <= 7'd0;
					9'b010110110: data_out <= 7'd0;
					9'b010110111: data_out <= 7'd0;
					9'b010111000: data_out <= 7'd0;
					9'b010111001: data_out <= 7'd0;
					9'b010111010: data_out <= 7'd0;
					9'b010111011: data_out <= 7'd0;
					9'b010111100: data_out <= 7'd0;
					9'b010111101: data_out <= 7'd0;
					9'b010111110: data_out <= 7'd0;
					9'b010111111: data_out <= 7'd0;
					9'b011000000: data_out <= 7'd0;
					9'b011000001: data_out <= 7'd0;
					9'b011000010: data_out <= 7'd0;
					9'b011000011: data_out <= 7'd0;
					9'b011000100: data_out <= 7'd0;
					9'b011000101: data_out <= 7'd0;
					9'b011000110: data_out <= 7'd0;
					9'b011000111: data_out <= 7'd0;
					9'b011001000: data_out <= 7'd0;
					9'b011001001: data_out <= 7'd0;
					9'b011001010: data_out <= 7'd0;
					9'b011001011: data_out <= 7'd0;
					9'b011001100: data_out <= 7'd0;
					9'b011001101: data_out <= 7'd0;
					9'b011001110: data_out <= 7'd0;
					9'b011001111: data_out <= 7'd0;
					9'b011010000: data_out <= 7'd0;
					9'b011010001: data_out <= 7'd0;
					9'b011010010: data_out <= 7'd0;
					9'b011010011: data_out <= 7'd0;
					9'b011010100: data_out <= 7'd0;
					9'b011010101: data_out <= 7'd0;
					9'b011010110: data_out <= 7'd0;
					9'b011010111: data_out <= 7'd0;
					9'b011011000: data_out <= 7'd0;
					9'b011011001: data_out <= 7'd0;
					9'b011011010: data_out <= 7'd0;
					9'b011011011: data_out <= 7'd0;
					9'b011011100: data_out <= 7'd0;
					9'b011011101: data_out <= 7'd0;
					9'b011011110: data_out <= 7'd0;
					9'b011011111: data_out <= 7'd0;
					9'b011100000: data_out <= 7'd0;
					9'b011100001: data_out <= 7'd0;
					9'b011100010: data_out <= 7'd0;
					9'b011100011: data_out <= 7'd0;
					9'b011100100: data_out <= 7'd0;
					9'b011100101: data_out <= 7'd0;
					9'b011100110: data_out <= 7'd0;
					9'b011100111: data_out <= 7'd0;
					9'b011101000: data_out <= 7'd0;
					9'b011101001: data_out <= 7'd0;
					9'b011101010: data_out <= 7'd0;
					9'b011101011: data_out <= 7'd0;
					9'b011101100: data_out <= 7'd0;
					9'b011101101: data_out <= 7'd0;
					9'b011101110: data_out <= 7'd0;
					9'b011101111: data_out <= 7'd0;
					9'b011110000: data_out <= 7'd0;
					9'b011110001: data_out <= 7'd0;
					9'b011110010: data_out <= 7'd0;
					9'b011110011: data_out <= 7'd0;
					9'b011110100: data_out <= 7'd0;
					9'b011110101: data_out <= 7'd0;
					9'b011110110: data_out <= 7'd0;
					9'b011110111: data_out <= 7'd0;
					9'b011111000: data_out <= 7'd0;
					9'b011111001: data_out <= 7'd0;
					9'b011111010: data_out <= 7'd0;
					9'b011111011: data_out <= 7'd0;
					9'b011111100: data_out <= 7'd0;
					9'b011111101: data_out <= 7'd0;
					9'b011111110: data_out <= 7'd0;
					9'b011111111: data_out <= 7'd0;
					9'b100000000: data_out <= 7'd2;
					9'b100000001: data_out <= 7'd2;
					9'b100000010: data_out <= 7'd4;
					9'b100000011: data_out <= 7'd4;
					9'b100000100: data_out <= 7'd2;
					9'b100000101: data_out <= 7'd2;
					9'b100000110: data_out <= 7'd6;
					9'b100000111: data_out <= 7'd7;
					9'b100001000: data_out <= 7'd8;
					9'b100001001: data_out <= 7'd4;
					9'b100001010: data_out <= 7'd4;
					9'b100001011: data_out <= 7'd10;
					9'b100001100: data_out <= 7'd12;
					9'b100001101: data_out <= 7'd16;
					9'b100001110: data_out <= 7'd19;
					9'b100001111: data_out <= 7'd20;
					9'b100010000: data_out <= 7'd21;
					9'b100010001: data_out <= 7'd12;
					9'b100010010: data_out <= 7'd22;
					9'b100010011: data_out <= 7'd23;
					9'b100010100: data_out <= 7'd24;
					9'b100010101: data_out <= 7'd25;
					9'b100010110: data_out <= 7'd30;
					9'b100010111: data_out <= 7'd31;
					9'b100011000: data_out <= 7'd32;
					9'b100011001: data_out <= 7'd33;
					9'b100011010: data_out <= 7'd34;
					9'b100011011: data_out <= 7'd35;
					9'b100011100: data_out <= 7'd36;
					9'b100011101: data_out <= 7'd37;
					9'b100011110: data_out <= 7'd39;
					9'b100011111: data_out <= 7'd41;
					9'b100100000: data_out <= 7'd42;
					9'b100100001: data_out <= 7'd43;
					9'b100100010: data_out <= 7'd44;
					9'b100100011: data_out <= 7'd45;
					9'b100100100: data_out <= 7'd46;
					9'b100100101: data_out <= 7'd48;
					9'b100100110: data_out <= 7'd49;
					9'b100100111: data_out <= 7'd50;
					9'b100101000: data_out <= 7'd51;
					9'b100101001: data_out <= 7'd52;
					9'b100101010: data_out <= 7'd53;
					9'b100101011: data_out <= 7'd54;
					9'b100101100: data_out <= 7'd55;
					9'b100101101: data_out <= 7'd56;
					9'b100101110: data_out <= 7'd43;
					9'b100101111: data_out <= 7'd44;
					9'b100110000: data_out <= 7'd45;
					9'b100110001: data_out <= 7'd58;
					9'b100110010: data_out <= 7'd59;
					9'b100110011: data_out <= 7'd60;
					9'b100110100: data_out <= 7'd61;
					9'b100110101: data_out <= 7'd62;
					9'b100110110: data_out <= 7'd3;
					9'b100110111: data_out <= 7'd61;
					9'b100111000: data_out <= 7'd62;
					9'b100111001: data_out <= 7'd63;
					9'b100111010: data_out <= 7'd64;
					9'b100111011: data_out <= 7'd62;
					9'b100111100: data_out <= 7'd65;
					9'b100111101: data_out <= 7'd3;
					9'b100111110: data_out <= 7'd64;
					9'b100111111: data_out <= 7'd62;
					9'b101000000: data_out <= 7'd66;

                    default: data_out = -1;

                endcase
            end
        
    endmodule